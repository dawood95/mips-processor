/*
  Everett Berry
  epberry@purdue.edu

  program counter
*/

`include "cpu_types_pkg.vh"

`include "datapath_cache_if.vh"

module pc (
  input logic CLK, nRST,
  datapath_cache_if.dp dpif
);

  //

endmodule
